scp Results.csv mihirm@ssh.pythonanywhere.com:valuemealstocks/
ssh mihirm@ssh.pythonanywhere.com
